module uart_tx(
	input x,
	output y
	);	

	assign y = x;
	
endmodule 