module rs232 (input x, output y);
	assign y = x;
endmodule 